module schematic-counter();

endmodule